`default_nettype none

module Task3
    (input logic start_game, grade_it, load_color,
     input logic [2:0] color_to_load,
     input logic [1:0] color_location,
     input logic [11:0] guess,
     output logic neopixel_data,
     output logic [3:0] round_number,
     output logic won, lost,
     input  logic clock, reset);




endmodule : Task3
